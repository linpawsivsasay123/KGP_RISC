`timescale 1ns / 1ps

module Diff_Module(Input, Output, Equal); 
    input [31:0] Input;
    output reg [31:0] Output; 
    output reg Equal; 

    wire [31:0] InputMinus1; 
    assign InputMinus1 = Input - 1;

    wire [31:0] InputMinus1XORInput; 
    wire [31:0] InputAndInputMinus1XORInput; 

    assign InputMinus1XORInput = InputMinus1 ^ Input; 
    assign InputAndInputMinus1XORInput = Input & InputMinus1XORInput;

    always @(*) begin
        case(InputAndInputMinus1XORInput)
            32'b00000000000000000000000000000001 : Output <= 0;
            32'b00000000000000000000000000000010 : Output <= 1;
            32'b00000000000000000000000000000100 : Output <= 2;
            32'b00000000000000000000000000001000 : Output <= 3;
            32'b00000000000000000000000000010000 : Output <= 4;
            32'b00000000000000000000000000100000 : Output <= 5;
            32'b00000000000000000000000001000000 : Output <= 6;
            32'b00000000000000000000000010000000 : Output <= 7;
            32'b00000000000000000000000100000000 : Output <= 8;
            32'b00000000000000000000001000000000 : Output <= 9;
            32'b00000000000000000000010000000000 : Output <= 10;
            32'b00000000000000000000100000000000 : Output <= 11;
            32'b00000000000000000001000000000000 : Output <= 12;
            32'b00000000000000000010000000000000 : Output <= 13;
            32'b00000000000000000100000000000000 : Output <= 14;
            32'b00000000000000001000000000000000 : Output <= 15;
            32'b00000000000000010000000000000000 : Output <= 16;
            32'b00000000000000100000000000000000 : Output <= 17;
            32'b00000000000001000000000000000000 : Output <= 18;
            32'b00000000000010000000000000000000 : Output <= 19;
            32'b00000000000100000000000000000000 : Output <= 20;
            32'b00000000001000000000000000000000 : Output <= 21;
            32'b00000000010000000000000000000000 : Output <= 22;
            32'b00000000100000000000000000000000 : Output <= 23;
            32'b00000001000000000000000000000000 : Output <= 24;
            32'b00000010000000000000000000000000 : Output <= 25;
            32'b00000100000000000000000000000000 : Output <= 26;
            32'b00001000000000000000000000000000 : Output <= 27;
            32'b00010000000000000000000000000000 : Output <= 28;
            32'b00100000000000000000000000000000 : Output <= 29;
            32'b01000000000000000000000000000000 : Output <= 30;
            32'b10000000000000000000000000000000 : Output <= 31;
        endcase
        if (InputAndInputMinus1XORInput == 32'd0)
            Equal <= 1;
        else
            Equal <= 0;
    end

endmodule